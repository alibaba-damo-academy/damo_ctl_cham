//////////////////////////////////////////////////
// Engineer: Chen Zhaohui (xinming)
// Email: chenzhaohui.czh@alibaba-inc.com
//
// Project Name: MVP
// Module Name: ntt_intt_defines
// Modify Date: 07/28/2021 11:10

// Description: Define timescale and some common params
//////////////////////////////////////////////////

`include "common_defines.vh"
`ifndef __NTT_INTT_DEFINES_VH__
`define __NTT_INTT_DEFINES_VH__

`define N 4096
`define  Q0 17314086913    // Q35 0
`define  Q1 17180393473    // Q35 1
`define  Q2 274886295553  // Q39

`endif // __NTT_INTT_DEFINES_VH__